(* tamara_triplicate *)
module top
#(parameter param291 = (((^~((&(8'hbd)) * ((8'hbd) <= (8'hb5)))) > (({(8'h9d), (8'ha3)} | (~^(8'hbe))) <<< {((8'hb0) ^ (7'h41))})) ? {(~|({(8'hb2), (8'h9f)} ? ((8'haa) ? (7'h42) : (8'hbc)) : (&(8'hb8)))), (({(8'hb1)} <<< (8'h9d)) >>> (((8'ha7) <<< (8'ha9)) ? (~|(8'hba)) : (8'h9d)))} : {{{((8'h9f) ? (8'hb7) : (8'hb5)), (&(8'hb1))}}, ({(~&(8'ha2)), {(8'hba)}} == (+{(8'h9f), (8'had)}))}),
parameter param292 = (|param291))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h14d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire0;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire signed [(5'h12):(1'h0)] wire2;
  input wire [(3'h4):(1'h0)] wire3;
  input wire [(2'h3):(1'h0)] wire4;
  wire signed [(3'h5):(1'h0)] wire289;
  wire [(4'hc):(1'h0)] wire288;
  wire signed [(2'h2):(1'h0)] wire287;
  wire [(3'h7):(1'h0)] wire286;
  wire [(5'h13):(1'h0)] wire284;
  wire [(5'h14):(1'h0)] wire279;
  wire signed [(5'h10):(1'h0)] wire278;
  wire [(4'hf):(1'h0)] wire277;
  wire signed [(4'he):(1'h0)] wire5;
  wire [(4'he):(1'h0)] wire6;
  wire [(5'h14):(1'h0)] wire7;
  wire signed [(5'h15):(1'h0)] wire8;
  wire signed [(4'hd):(1'h0)] wire9;
  wire [(5'h11):(1'h0)] wire10;
  wire signed [(5'h14):(1'h0)] wire11;
  wire signed [(2'h2):(1'h0)] wire12;
  wire signed [(5'h12):(1'h0)] wire13;
  wire [(5'h15):(1'h0)] wire14;
  wire signed [(3'h6):(1'h0)] wire15;
  wire [(4'hf):(1'h0)] wire275;
  reg [(5'h15):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg281 = (1'h0);
  assign y = {wire289,
                 wire288,
                 wire287,
                 wire286,
                 wire284,
                 wire279,
                 wire278,
                 wire277,
                 wire5,
                 wire6,
                 wire7,
                 wire8,
                 wire9,
                 wire10,
                 wire11,
                 wire12,
                 wire13,
                 wire14,
                 wire15,
                 wire275,
                 reg283,
                 reg282,
                 reg281,
                 (1'h0)};
  assign wire5 = $unsigned((^~wire0[(3'h4):(3'h4)]));
  assign wire6 = (8'had);
  assign wire7 = wire2[(1'h0):(1'h0)];
  assign wire8 = wire3;
  assign wire9 = wire0;
  assign wire10 = (|wire9[(3'h7):(2'h2)]);
  assign wire11 = wire3[(2'h2):(1'h0)];
  assign wire12 = wire7[(4'hb):(4'ha)];
  assign wire13 = $unsigned((^(^$signed(wire5))));
  assign wire14 = wire7[(4'hd):(2'h3)];
  assign wire15 = (^wire12);
  module16 #() modinst276 (wire275, clk, wire13, wire0, wire5, wire7, wire14);
  assign wire277 = (($unsigned(($signed(wire14) ?
                           $unsigned(wire9) : $unsigned(wire275))) || $unsigned({(wire5 ?
                               wire275 : wire15),
                           $signed(wire9)})) ?
                       ({((8'had) ?
                               wire14 : $signed(wire0))} || $signed(wire9)) : wire5[(2'h2):(1'h1)]);
  assign wire278 = wire13[(4'ha):(4'ha)];
  module111 #() modinst280 (wire279, clk, wire6, wire15, wire14, wire278);
  always
    @(posedge clk) begin
      reg281 <= $signed((wire4[(2'h2):(2'h2)] || ({(&wire12),
          $unsigned(wire279)} << wire4[(1'h1):(1'h1)])));
      reg282 <= $signed({wire4});
      reg283 <= (^(({((8'ha3) ? (8'hb2) : wire7),
          $unsigned(wire10)} >>> $unsigned((wire4 ?
          wire11 : wire7))) ~^ $signed({(~|wire278), (wire15 | wire6)})));
    end
  module111 #() modinst285 (wire284, clk, wire14, wire7, wire277, wire1);
  assign wire286 = $signed($unsigned((~^$unsigned(wire10))));
  assign wire287 = wire286;
  assign wire288 = wire277;
  module173 #() modinst290 (.wire174(wire284), .y(wire289), .wire177(wire11), .clk(clk), .wire176(wire13), .wire175(wire277));
endmodule

module module16
#(parameter param273 = ((8'hbb) ? (((~(~^(8'hb1))) ? ({(8'hbf)} ? {(8'hba)} : (7'h44)) : ((+(7'h42)) | (+(8'hbd)))) ? (8'hb5) : ({{(8'hbc)}} ? (^~(&(8'hba))) : (8'hbe))) : {((((8'hbf) < (8'ha7)) <= (-(8'ha8))) ? ((!(7'h43)) ? ((8'ha1) < (8'h9c)) : (|(8'h9f))) : {((8'hbf) ? (8'ha3) : (8'hae)), (~^(8'hbe))})}),
parameter param274 = (!(({(param273 ? param273 : param273)} ~^ {(^~param273)}) | param273)))
(y, clk, wire17, wire18, wire19, wire20, wire21);
  output wire [(32'h1fb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire17;
  input wire [(5'h14):(1'h0)] wire18;
  input wire [(4'he):(1'h0)] wire19;
  input wire [(5'h14):(1'h0)] wire20;
  input wire [(4'he):(1'h0)] wire21;
  wire [(4'ha):(1'h0)] wire22;
  wire signed [(3'h6):(1'h0)] wire74;
  wire [(5'h15):(1'h0)] wire76;
  wire signed [(5'h11):(1'h0)] wire77;
  wire signed [(2'h2):(1'h0)] wire102;
  wire signed [(5'h11):(1'h0)] wire104;
  wire signed [(4'h9):(1'h0)] wire105;
  wire [(4'hf):(1'h0)] wire106;
  wire signed [(5'h15):(1'h0)] wire107;
  wire signed [(3'h4):(1'h0)] wire108;
  wire [(5'h15):(1'h0)] wire109;
  wire signed [(4'hf):(1'h0)] wire110;
  wire [(5'h13):(1'h0)] wire162;
  wire [(2'h2):(1'h0)] wire164;
  wire signed [(4'ha):(1'h0)] wire210;
  wire [(4'hb):(1'h0)] wire212;
  wire [(5'h11):(1'h0)] wire227;
  wire signed [(2'h3):(1'h0)] wire271;
  reg signed [(4'hf):(1'h0)] reg226 = (1'h0);
  reg [(4'h8):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg222 = (1'h0);
  reg [(3'h7):(1'h0)] reg221 = (1'h0);
  reg [(4'hd):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg219 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg217 = (1'h0);
  reg [(5'h13):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg215 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg214 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg213 = (1'h0);
  reg [(5'h15):(1'h0)] reg172 = (1'h0);
  reg [(4'ha):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg167 = (1'h0);
  reg [(4'hf):(1'h0)] reg166 = (1'h0);
  reg [(4'ha):(1'h0)] reg165 = (1'h0);
  assign y = {wire22,
                 wire74,
                 wire76,
                 wire77,
                 wire102,
                 wire104,
                 wire105,
                 wire106,
                 wire107,
                 wire108,
                 wire109,
                 wire110,
                 wire162,
                 wire164,
                 wire210,
                 wire212,
                 wire227,
                 wire271,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 (1'h0)};
  assign wire22 = wire21;
  module23 #() modinst75 (.wire25(wire20), .y(wire74), .wire24(wire17), .clk(clk), .wire26(wire18), .wire27(wire22));
  assign wire76 = $signed((-($unsigned($unsigned(wire17)) ?
                      ({wire20, wire20} ?
                          {wire74, wire20} : wire22) : $signed((wire17 ?
                          wire74 : wire20)))));
  assign wire77 = (wire76 ?
                      wire20 : (wire74 ?
                          (~&$unsigned({wire17})) : (wire21 ?
                              $unsigned($unsigned(wire76)) : ((wire20 ?
                                  wire74 : wire19) | wire18))));
  module78 #() modinst103 (.wire82(wire19), .wire80(wire77), .wire81(wire76), .clk(clk), .wire79(wire20), .y(wire102));
  assign wire104 = ((wire22[(3'h5):(3'h4)] <<< $unsigned((wire77[(4'hc):(4'hb)] ^~ wire19))) ?
                       {wire102[(1'h1):(1'h1)],
                           $signed({wire77[(4'h8):(2'h3)]})} : $signed((^(-(wire76 && wire21)))));
  assign wire105 = $signed((!(!(wire76 || (&wire22)))));
  assign wire106 = $unsigned(wire74[(3'h4):(1'h1)]);
  assign wire107 = wire104;
  assign wire108 = ($unsigned((|($signed(wire20) ?
                           wire19[(3'h4):(2'h2)] : $unsigned(wire77)))) ?
                       (^wire22[(3'h4):(1'h1)]) : $unsigned(wire20));
  assign wire109 = wire102[(2'h2):(1'h0)];
  assign wire110 = (-$unsigned({((wire105 ? (8'hbc) : wire108) ?
                           $signed(wire107) : $unsigned(wire21)),
                       $unsigned(((8'ha4) >>> wire22))}));
  module111 #() modinst163 (.wire115(wire19), .wire114(wire102), .y(wire162), .wire113(wire21), .wire112(wire18), .clk(clk));
  assign wire164 = (8'hac);
  always
    @(posedge clk) begin
      reg165 <= $signed(wire104);
      reg166 <= $unsigned($signed(wire164[(2'h2):(1'h1)]));
      reg167 <= wire104;
      if ((^((((wire110 ? wire22 : wire106) ?
              $signed(wire105) : $unsigned(wire76)) ?
          $unsigned((reg167 ?
              wire105 : wire162)) : ($unsigned(reg165) >= (wire19 ?
              wire107 : wire108))) + reg167[(1'h0):(1'h0)])))
        begin
          reg168 <= (wire19[(4'h8):(3'h6)] || $signed(wire19[(3'h5):(3'h4)]));
          reg169 <= wire18[(5'h10):(4'hd)];
          reg170 <= wire109[(3'h4):(2'h2)];
          reg171 <= (wire104 << (8'hb5));
        end
      else
        begin
          reg168 <= {wire19, wire74[(1'h0):(1'h0)]};
          reg169 <= ((8'h9e) == (8'ha5));
        end
      reg172 <= (~(reg167 ? wire110[(1'h1):(1'h1)] : reg170[(4'hb):(3'h4)]));
    end
  module173 #() modinst211 (wire210, clk, wire20, reg170, reg166, wire109);
  assign wire212 = (&{reg171[(2'h3):(2'h3)]});
  always
    @(posedge clk) begin
      if (wire74[(2'h2):(1'h1)])
        begin
          reg213 <= $signed({reg166});
          if ($unsigned(reg166))
            begin
              reg214 <= (~|wire108);
              reg215 <= ($unsigned((~wire74)) ^ (($signed((^~wire19)) ?
                  $unsigned((wire108 || (8'hae))) : $unsigned((wire106 ?
                      wire20 : wire102))) >>> ($signed((wire74 ?
                  wire162 : wire110)) <= (reg170 ?
                  (wire106 ? wire105 : reg171) : (wire106 & reg170)))));
              reg216 <= (($unsigned(reg166) ?
                  $signed(((wire74 ? (8'hb8) : (7'h43)) ?
                      wire22 : $signed(reg165))) : (((~&wire108) ?
                          $signed(wire77) : (reg168 ? (8'ha1) : wire109)) ?
                      wire162[(4'hc):(3'h5)] : reg166[(4'ha):(3'h5)])) <= wire106);
              reg217 <= (({$signed($signed(reg171)), wire212[(3'h7):(3'h4)]} ?
                      (wire77[(1'h0):(1'h0)] ?
                          ({reg169, wire162} ?
                              reg169 : reg169) : $signed((reg213 ?
                              wire162 : wire210))) : (!$signed((wire104 + reg169)))) ?
                  wire74[(2'h3):(2'h2)] : (((+(-wire18)) >> $unsigned((+wire164))) < wire21[(4'h9):(2'h3)]));
            end
          else
            begin
              reg214 <= $signed(wire76[(1'h0):(1'h0)]);
            end
          reg218 <= wire17;
        end
      else
        begin
          if (wire106)
            begin
              reg213 <= (($signed({wire104[(3'h7):(2'h2)]}) && (~|($signed(reg214) >> (reg213 ?
                  wire104 : reg172)))) <= $signed((~|wire210)));
              reg214 <= {reg214[(2'h2):(2'h2)]};
            end
          else
            begin
              reg213 <= $signed(((wire212[(3'h7):(3'h4)] * ((wire105 || reg165) ?
                  (8'ha7) : {wire74, wire109})) && wire102));
              reg214 <= ($signed(reg166[(4'hb):(2'h3)]) ?
                  $unsigned($signed({$signed((8'hab)), (^wire76)})) : wire21);
              reg215 <= (~$unsigned((($signed(wire162) ^~ $signed(reg214)) ?
                  ($signed(reg172) ?
                      (reg172 ? (8'haf) : wire18) : (reg167 ?
                          reg218 : wire76)) : wire164[(2'h2):(1'h1)])));
              reg216 <= (^~(^~reg168[(1'h0):(1'h0)]));
              reg217 <= (wire109[(3'h4):(1'h0)] ?
                  ((~|wire104[(4'h9):(3'h7)]) ?
                      $unsigned((^~wire164)) : ({(reg214 ? reg167 : wire106),
                          $signed((8'hb0))} <<< {$signed(wire212)})) : wire108[(1'h1):(1'h0)]);
            end
        end
      if ((~(!$unsigned(wire19))))
        begin
          reg219 <= $signed($signed(reg215));
          reg220 <= (~$unsigned((((reg218 ? wire18 : wire17) ?
                  (wire105 ? (8'hb3) : wire210) : wire76) ?
              (reg218 + (wire162 ? wire212 : reg215)) : reg171)));
          reg221 <= {(wire212 ?
                  ($unsigned(reg165[(1'h1):(1'h1)]) != reg220) : $signed($unsigned((+reg217)))),
              ((|{reg169}) ?
                  (+$unsigned((reg172 ?
                      wire110 : wire107))) : ($signed((^~reg220)) - reg214[(2'h2):(1'h0)]))};
          reg222 <= $unsigned($unsigned(wire21));
        end
      else
        begin
          reg219 <= ((-$signed((reg169 ? (reg222 > wire76) : wire17))) ?
              $unsigned((~&(8'ha5))) : wire18[(1'h1):(1'h1)]);
          if ($signed(reg221))
            begin
              reg220 <= $signed($unsigned(($unsigned((reg218 > reg222)) ?
                  (wire74 ?
                      (reg214 ?
                          wire108 : reg221) : wire20) : $unsigned(wire104[(5'h11):(4'h9)]))));
              reg221 <= (~^{($signed($unsigned(reg218)) | $signed(wire20)),
                  (|{$unsigned(reg221), $unsigned(reg167)})});
              reg222 <= wire19;
              reg223 <= (reg220 && reg169[(1'h1):(1'h0)]);
              reg224 <= $unsigned(wire109[(4'ha):(3'h4)]);
            end
          else
            begin
              reg220 <= (($signed((wire162[(3'h7):(3'h5)] ?
                  $signed(wire105) : (8'hb9))) || (wire22[(4'h9):(1'h1)] >>> $signed((+reg219)))) + (wire212[(1'h0):(1'h0)] ?
                  $unsigned($unsigned((7'h42))) : $unsigned(reg165)));
            end
          reg225 <= $signed(((^~((8'hb3) ?
              $signed(reg218) : (8'hb1))) * (8'h9e)));
        end
      reg226 <= $signed(reg216);
    end
  assign wire227 = $unsigned($signed($signed(($signed((8'hac)) ^~ wire17[(1'h0):(1'h0)]))));
  module228 #() modinst272 (.wire232(wire76), .wire231(reg169), .wire233(reg213), .y(wire271), .clk(clk), .wire229(wire227), .wire230(wire105));
endmodule

module module228
#(parameter param269 = ((((!{(7'h42), (8'hb8)}) ? (((8'hb0) ? (8'ha8) : (7'h41)) ? ((8'hb6) >> (8'ha3)) : ((8'ha7) ? (7'h44) : (8'haf))) : ((8'ha5) * (^(8'ha1)))) < ((((8'hb0) >= (8'hbb)) ? ((8'hbf) || (8'ha5)) : ((8'hb8) ? (8'hac) : (8'ha9))) * ((|(7'h42)) << {(8'h9e), (7'h44)}))) ? (^((8'ha6) | (((8'ha5) ~^ (7'h40)) ? (!(8'hba)) : (~|(8'ha4))))) : (((((8'hbd) <<< (8'ha6)) ? ((8'hab) != (8'hac)) : ((8'hb5) ~^ (8'hbf))) ? (7'h43) : (((8'h9e) + (8'ha5)) ? {(8'h9d)} : {(8'ha0), (8'hb1)})) << (((!(8'hb6)) != (~^(8'hb0))) < (((8'h9e) ? (8'hbf) : (8'hb5)) > ((8'hbc) ? (8'hb8) : (8'ha2)))))),
parameter param270 = (param269 ? (((-(+param269)) ? (((8'ha3) >>> param269) ? ((8'haa) ? param269 : param269) : param269) : param269) >> (param269 >> {(param269 ^~ param269)})) : param269))
(y, clk, wire233, wire232, wire231, wire230, wire229);
  output wire [(32'h1a4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire233;
  input wire signed [(5'h11):(1'h0)] wire232;
  input wire signed [(5'h13):(1'h0)] wire231;
  input wire [(3'h4):(1'h0)] wire230;
  input wire signed [(5'h11):(1'h0)] wire229;
  wire [(5'h11):(1'h0)] wire268;
  wire [(4'hb):(1'h0)] wire255;
  wire [(4'hc):(1'h0)] wire254;
  wire [(4'hd):(1'h0)] wire253;
  wire signed [(3'h4):(1'h0)] wire252;
  wire [(4'hd):(1'h0)] wire250;
  wire [(5'h11):(1'h0)] wire249;
  wire signed [(5'h14):(1'h0)] wire243;
  wire signed [(4'h8):(1'h0)] wire241;
  wire [(3'h6):(1'h0)] wire240;
  wire signed [(5'h10):(1'h0)] wire239;
  wire signed [(5'h11):(1'h0)] wire238;
  reg signed [(3'h6):(1'h0)] reg267 = (1'h0);
  reg [(4'hf):(1'h0)] reg266 = (1'h0);
  reg [(5'h13):(1'h0)] reg265 = (1'h0);
  reg [(4'hb):(1'h0)] reg264 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg263 = (1'h0);
  reg [(4'he):(1'h0)] reg262 = (1'h0);
  reg signed [(4'he):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg260 = (1'h0);
  reg [(5'h12):(1'h0)] reg259 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg258 = (1'h0);
  reg [(4'hf):(1'h0)] reg257 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg256 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg247 = (1'h0);
  reg [(4'h9):(1'h0)] reg246 = (1'h0);
  reg [(4'hc):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg244 = (1'h0);
  reg [(5'h15):(1'h0)] reg242 = (1'h0);
  reg [(4'he):(1'h0)] reg237 = (1'h0);
  reg [(3'h6):(1'h0)] reg236 = (1'h0);
  reg [(4'h8):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg234 = (1'h0);
  assign y = {wire268,
                 wire255,
                 wire254,
                 wire253,
                 wire252,
                 wire250,
                 wire249,
                 wire243,
                 wire241,
                 wire240,
                 wire239,
                 wire238,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg251,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg242,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed((wire232 ? (&$unsigned({wire232})) : (8'hbd))))
        begin
          reg234 <= $unsigned((|(-wire230)));
        end
      else
        begin
          reg234 <= wire232;
        end
      reg235 <= ((-$signed(wire231[(3'h5):(3'h4)])) || ($unsigned(wire230) ?
          (&wire232[(4'hc):(1'h0)]) : (((+wire232) ?
              (wire233 ?
                  wire231 : (8'ha5)) : $unsigned(wire229)) << (~^(wire229 ~^ reg234)))));
      reg236 <= wire229;
      reg237 <= (reg235[(1'h0):(1'h0)] ?
          ((-(~|(wire231 ? wire233 : reg235))) ?
              ((+$unsigned(wire231)) ?
                  $unsigned((wire229 ?
                      (8'hba) : wire230)) : wire229) : $unsigned((wire230[(3'h4):(3'h4)] < (reg236 ?
                  (8'ha2) : wire233)))) : (|{(~|(reg236 ? reg236 : reg234)),
              $signed(reg236)}));
    end
  assign wire238 = {(($signed((!reg234)) ~^ reg236) ?
                           $signed(wire230) : (~&(|wire231[(4'h9):(1'h1)]))),
                       wire231[(4'h9):(2'h3)]};
  assign wire239 = reg236;
  assign wire240 = wire230[(2'h2):(2'h2)];
  assign wire241 = wire240[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg242 <= (-wire231);
    end
  assign wire243 = $signed(((+$unsigned((reg237 ^ wire240))) ?
                       wire241 : $unsigned(wire232)));
  always
    @(posedge clk) begin
      reg244 <= reg234[(3'h6):(3'h6)];
      reg245 <= $signed(wire231[(4'hb):(1'h1)]);
      if ((+$unsigned(($signed((wire233 != wire232)) ?
          (&$unsigned(wire230)) : wire232[(1'h0):(1'h0)]))))
        begin
          reg246 <= (reg242 ?
              $signed((^((-wire233) == $signed(wire229)))) : ($unsigned(reg235) ?
                  (~|((~reg236) ?
                      (~|reg234) : wire229[(3'h4):(1'h0)])) : $signed(reg244)));
          reg247 <= wire231;
        end
      else
        begin
          reg246 <= (|($unsigned(wire243) & (^{wire232[(4'hb):(4'hb)],
              (reg244 ? reg237 : (7'h40))})));
          reg247 <= wire233[(4'h8):(3'h6)];
          reg248 <= $unsigned($unsigned(reg246[(1'h0):(1'h0)]));
        end
    end
  assign wire249 = $signed((((~&reg242[(4'hc):(4'ha)]) & (~^$unsigned(wire229))) << reg247));
  assign wire250 = ($unsigned(($signed((~&wire249)) ?
                           reg234[(4'h9):(3'h4)] : $signed((^wire243)))) ?
                       $signed($unsigned((wire233 ^ ((8'hb1) ?
                           wire238 : reg248)))) : $unsigned(reg245));
  always
    @(posedge clk) begin
      reg251 <= $unsigned({reg242,
          {($unsigned(reg247) >= (^~wire230)),
              ({reg247, reg242} ? $unsigned((8'hbc)) : (~&wire239))}});
    end
  assign wire252 = $signed((^~({{reg236}} >>> $unsigned($unsigned(wire239)))));
  assign wire253 = ($signed((8'hbb)) != $signed($unsigned((!$signed(wire232)))));
  assign wire254 = ((reg247 ?
                           wire240[(2'h2):(1'h1)] : ((~|$unsigned(wire253)) ?
                               wire231[(2'h3):(2'h3)] : reg245[(1'h1):(1'h1)])) ?
                       (!(reg245 ?
                           (wire231 ?
                               (~&reg246) : (wire233 ^ reg242)) : (((8'ha3) ?
                                   wire253 : wire240) ?
                               $unsigned(wire232) : $unsigned(wire243)))) : ($unsigned(($unsigned(wire249) & $signed((7'h44)))) | ($signed((+(8'ha8))) ~^ $signed((reg237 == wire252)))));
  assign wire255 = (^wire250[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg256 <= reg235[(1'h0):(1'h0)];
      reg257 <= ($signed(wire252[(1'h1):(1'h0)]) ?
          reg235 : wire255[(4'hb):(4'ha)]);
      if (($signed({{(wire243 ? reg235 : reg237)}}) | wire231))
        begin
          reg258 <= (((~^reg234[(2'h2):(2'h2)]) ?
                  $unsigned({(wire241 ^~ wire231),
                      {reg256, reg242}}) : $unsigned(((reg237 ?
                          wire230 : wire233) ?
                      $signed(reg256) : (wire255 && wire238)))) ?
              reg248 : $unsigned((^~wire233)));
          reg259 <= $signed({$signed($signed($unsigned(wire253)))});
          reg260 <= wire252[(1'h0):(1'h0)];
          if (((!reg242) <= $unsigned($signed((wire241[(1'h1):(1'h1)] & {wire231})))))
            begin
              reg261 <= reg247[(3'h6):(2'h2)];
            end
          else
            begin
              reg261 <= reg260;
              reg262 <= {(8'hb7),
                  ($unsigned(wire255) ?
                      $unsigned(((^~wire254) ?
                          $signed(wire233) : {reg251})) : {wire253})};
              reg263 <= wire230;
              reg264 <= $unsigned(({((wire233 ? wire241 : reg261) ?
                          {reg242, reg246} : $signed(wire253))} ?
                  wire253 : reg251[(1'h0):(1'h0)]));
            end
        end
      else
        begin
          reg258 <= reg256[(2'h2):(2'h2)];
          reg259 <= {$unsigned(((~&reg244) ?
                  $unsigned((wire230 ? wire241 : wire254)) : reg264)),
              wire249};
          reg260 <= $unsigned((({$unsigned(wire250)} ?
                  ((reg256 ? wire232 : reg257) ?
                      (reg263 ?
                          wire243 : wire250) : (reg264 != reg251)) : $unsigned($unsigned(reg247))) ?
              {$unsigned($unsigned(wire233))} : {$unsigned($unsigned((8'hb4)))}));
        end
    end
  always
    @(posedge clk) begin
      reg265 <= $signed($unsigned(($unsigned((wire240 ? reg261 : (8'h9f))) ?
          (((8'hab) ? (8'hb6) : reg257) ?
              wire239 : reg259[(4'h9):(3'h5)]) : $unsigned((|wire230)))));
      reg266 <= {wire230[(2'h2):(2'h2)], {reg264[(4'h9):(3'h6)]}};
    end
  always
    @(posedge clk) begin
      reg267 <= wire254[(1'h1):(1'h1)];
    end
  assign wire268 = $unsigned({wire229});
endmodule

module module173  (y, clk, wire177, wire176, wire175, wire174);
  output wire [(32'h13e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire177;
  input wire signed [(5'h12):(1'h0)] wire176;
  input wire [(4'hf):(1'h0)] wire175;
  input wire signed [(4'hd):(1'h0)] wire174;
  wire signed [(5'h13):(1'h0)] wire209;
  wire signed [(3'h6):(1'h0)] wire208;
  wire signed [(3'h5):(1'h0)] wire207;
  wire signed [(4'ha):(1'h0)] wire206;
  wire [(2'h3):(1'h0)] wire205;
  wire signed [(4'hd):(1'h0)] wire204;
  wire [(2'h3):(1'h0)] wire200;
  wire signed [(3'h7):(1'h0)] wire199;
  wire [(4'hc):(1'h0)] wire198;
  wire [(4'h9):(1'h0)] wire197;
  wire [(4'hb):(1'h0)] wire196;
  wire signed [(4'hb):(1'h0)] wire185;
  wire signed [(3'h7):(1'h0)] wire184;
  wire [(2'h2):(1'h0)] wire183;
  wire [(4'hd):(1'h0)] wire179;
  reg signed [(5'h10):(1'h0)] reg203 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg202 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg194 = (1'h0);
  reg [(2'h2):(1'h0)] reg193 = (1'h0);
  reg [(4'hb):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg191 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg190 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg189 = (1'h0);
  reg [(5'h13):(1'h0)] reg188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg186 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg [(5'h11):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg178 = (1'h0);
  assign y = {wire209,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 wire196,
                 wire185,
                 wire184,
                 wire183,
                 wire179,
                 reg203,
                 reg202,
                 reg201,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg182,
                 reg181,
                 reg180,
                 reg178,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg178 <= {(|$unsigned($unsigned(((8'had) ? wire177 : wire174))))};
    end
  assign wire179 = (wire175[(3'h5):(1'h1)] ? wire177 : reg178);
  always
    @(posedge clk) begin
      reg180 <= (($signed((wire179 || (wire177 < wire179))) <<< wire176) ?
          $signed($signed((wire176 ^ $unsigned(reg178)))) : ((reg178 & wire175[(1'h1):(1'h0)]) ?
              $signed($unsigned(wire179)) : $signed(reg178)));
      reg181 <= $unsigned({(+(~|$unsigned(reg180)))});
      reg182 <= reg181;
    end
  assign wire183 = {(reg180[(2'h3):(1'h0)] ?
                           (|(!$unsigned(wire177))) : $unsigned($signed(reg181))),
                       (|$signed($unsigned((8'hac))))};
  assign wire184 = (wire175[(4'hb):(3'h5)] ?
                       $unsigned((!reg182[(3'h5):(2'h3)])) : wire179[(3'h5):(1'h0)]);
  assign wire185 = wire177;
  always
    @(posedge clk) begin
      if ((-wire179[(2'h2):(2'h2)]))
        begin
          reg186 <= ((reg180 - (^~{(reg182 > wire176),
              {wire177,
                  wire177}})) <<< (wire175[(2'h2):(1'h0)] <<< (reg180 ~^ ($unsigned(wire179) ?
              {reg178, wire175} : $unsigned(wire185)))));
        end
      else
        begin
          reg186 <= {((+(^(wire185 >= reg180))) ?
                  wire174[(4'h8):(3'h7)] : (^~reg182))};
          reg187 <= ((($signed((^reg186)) ?
              {wire179, (wire183 ? wire185 : wire176)} : ((reg180 ?
                      wire174 : wire179) ?
                  {reg178,
                      wire179} : (~|wire179))) | $signed(((wire185 >>> reg178) ?
              (reg181 << wire184) : wire175[(4'hf):(3'h6)]))) >> wire174);
        end
      if ((wire177 ?
          (^~(~(reg181 ? {reg187} : (!reg178)))) : reg186[(3'h5):(3'h4)]))
        begin
          if ({wire176[(3'h6):(2'h2)]})
            begin
              reg188 <= ((wire183[(1'h0):(1'h0)] ?
                  (reg180 & $unsigned(reg178)) : ((wire177 >> (reg181 >> wire179)) ?
                      {reg180,
                          (reg181 ?
                              (8'ha5) : wire175)} : {(wire175 || wire174)})) < (~^$unsigned((~^reg181[(5'h11):(3'h4)]))));
            end
          else
            begin
              reg188 <= ({(^~({wire176, wire177} ?
                      (wire177 ^ wire179) : (reg181 >> wire184)))} & ($signed(reg186[(3'h7):(3'h4)]) ?
                  $signed(({wire174,
                      wire175} > (wire185 || wire174))) : $unsigned($signed($signed(wire179)))));
              reg189 <= reg182;
              reg190 <= (((reg188 & reg178[(3'h6):(1'h1)]) ?
                      wire185[(1'h0):(1'h0)] : $signed($signed(wire177))) ?
                  wire184 : reg182);
              reg191 <= reg186[(3'h5):(3'h5)];
              reg192 <= $signed(((($unsigned((8'hbf)) ? (8'hac) : (~&reg188)) ?
                      $signed((wire175 ?
                          (8'hb5) : reg187)) : reg186[(1'h1):(1'h1)]) ?
                  $signed(reg180) : $signed($unsigned($signed(reg191)))));
            end
          reg193 <= $unsigned(reg191);
          reg194 <= (&{(~|(^~reg190))});
          reg195 <= ((~&$signed({(reg194 ^ (8'hb5)), (8'hb3)})) | wire184);
        end
      else
        begin
          reg188 <= ({(~|($unsigned(reg182) | (wire185 == reg192)))} | reg191[(4'ha):(1'h1)]);
        end
    end
  assign wire196 = (~&wire185);
  assign wire197 = (8'hb2);
  assign wire198 = $unsigned(({reg188[(3'h4):(1'h0)]} ?
                       $signed(wire175) : $unsigned(reg188[(2'h3):(2'h3)])));
  assign wire199 = reg187[(4'h9):(3'h4)];
  assign wire200 = ((((|{wire185}) && ($unsigned(reg186) <= (reg187 * reg194))) << (({reg186,
                               reg193} ?
                           reg180[(2'h3):(1'h0)] : $signed((8'hbb))) < (~|wire175[(1'h0):(1'h0)]))) ?
                       {(-$unsigned($unsigned(wire177)))} : (|reg186));
  always
    @(posedge clk) begin
      reg201 <= $unsigned($unsigned($unsigned({(wire176 | wire176), wire185})));
      reg202 <= (wire183 ?
          $unsigned($unsigned((reg201 ?
              (^~reg192) : reg178))) : ($signed(wire175) + wire175));
      reg203 <= reg192;
    end
  assign wire204 = reg188[(4'ha):(3'h7)];
  assign wire205 = wire197;
  assign wire206 = (~^(({(!wire199), {(8'hba), wire175}} <<< (~&(wire174 ?
                           wire176 : wire199))) ?
                       $signed((|$signed(reg181))) : ({((8'ha2) != wire183)} << wire179[(4'hb):(3'h4)])));
  assign wire207 = (&(8'ha7));
  assign wire208 = $unsigned((reg203 || $unsigned({$signed((8'ha1)),
                       (wire196 ? reg187 : wire207)})));
  assign wire209 = reg182;
endmodule

module module111
#(parameter param161 = (((8'ha9) || (8'h9e)) << (((+((7'h44) ? (8'hb4) : (8'h9d))) <<< (&(~^(8'h9c)))) ? (~&(((8'hae) ? (8'hb4) : (8'h9f)) ? {(8'hb7), (8'hb9)} : ((7'h42) ? (8'ha5) : (8'hbb)))) : (~|(!{(8'ha0), (8'hb8)})))))
(y, clk, wire115, wire114, wire113, wire112);
  output wire [(32'h204):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire115;
  input wire signed [(2'h2):(1'h0)] wire114;
  input wire signed [(4'he):(1'h0)] wire113;
  input wire [(5'h10):(1'h0)] wire112;
  wire signed [(5'h14):(1'h0)] wire160;
  wire signed [(2'h3):(1'h0)] wire146;
  wire signed [(4'hc):(1'h0)] wire145;
  wire [(4'ha):(1'h0)] wire144;
  wire signed [(3'h4):(1'h0)] wire143;
  wire signed [(5'h12):(1'h0)] wire142;
  wire signed [(4'h9):(1'h0)] wire141;
  wire signed [(3'h6):(1'h0)] wire123;
  wire [(5'h13):(1'h0)] wire120;
  wire [(5'h14):(1'h0)] wire118;
  wire signed [(5'h13):(1'h0)] wire117;
  wire [(4'h9):(1'h0)] wire116;
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg157 = (1'h0);
  reg [(5'h10):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg153 = (1'h0);
  reg [(2'h3):(1'h0)] reg152 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg150 = (1'h0);
  reg [(5'h11):(1'h0)] reg149 = (1'h0);
  reg [(4'he):(1'h0)] reg148 = (1'h0);
  reg [(5'h14):(1'h0)] reg147 = (1'h0);
  reg [(4'ha):(1'h0)] reg140 = (1'h0);
  reg [(4'hf):(1'h0)] reg139 = (1'h0);
  reg [(5'h13):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg137 = (1'h0);
  reg [(4'h8):(1'h0)] reg136 = (1'h0);
  reg [(4'hd):(1'h0)] reg135 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg134 = (1'h0);
  reg [(4'h9):(1'h0)] reg133 = (1'h0);
  reg [(4'he):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg131 = (1'h0);
  reg [(3'h5):(1'h0)] reg130 = (1'h0);
  reg [(5'h13):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg127 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg125 = (1'h0);
  reg [(4'hb):(1'h0)] reg124 = (1'h0);
  reg [(5'h15):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg121 = (1'h0);
  reg [(5'h11):(1'h0)] reg119 = (1'h0);
  assign y = {wire160,
                 wire146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire123,
                 wire120,
                 wire118,
                 wire117,
                 wire116,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg122,
                 reg121,
                 reg119,
                 (1'h0)};
  assign wire116 = wire115;
  assign wire117 = $signed(wire115);
  assign wire118 = ({$signed($unsigned(wire113[(2'h3):(1'h0)])),
                       $signed((wire117 - (~^wire114)))} >> {(wire116 ?
                           wire112[(4'hf):(3'h6)] : ((wire115 ?
                                   wire112 : wire117) ?
                               $signed(wire113) : $unsigned(wire116))),
                       $signed((!wire114))});
  always
    @(posedge clk) begin
      reg119 <= wire115[(4'he):(1'h0)];
    end
  assign wire120 = wire118[(4'h8):(3'h6)];
  always
    @(posedge clk) begin
      reg121 <= (!wire114[(1'h1):(1'h0)]);
      reg122 <= $unsigned((+(((wire112 >>> (8'ha0)) >= (wire117 ?
          wire114 : (8'hbd))) != wire112[(2'h2):(1'h0)])));
    end
  assign wire123 = (wire118[(4'hc):(4'hb)] ?
                       (($signed({reg121, reg121}) ?
                           wire112 : $signed($signed(reg119))) != {$unsigned($signed(wire120)),
                           $unsigned(reg122[(5'h15):(3'h5)])}) : $unsigned(((reg121 ^ (wire120 >= wire113)) ?
                           (&(8'h9e)) : reg121[(2'h2):(1'h1)])));
  always
    @(posedge clk) begin
      if (reg122)
        begin
          reg124 <= $unsigned($unsigned($unsigned($signed($signed(wire112)))));
        end
      else
        begin
          if (($signed((+$signed((reg119 >> wire118)))) - {(-((~reg122) ^~ ((7'h42) ^~ wire113))),
              {reg119, $unsigned(wire113[(1'h0):(1'h0)])}}))
            begin
              reg124 <= ((&$signed({wire117[(1'h0):(1'h0)]})) * $unsigned($signed(($unsigned((8'hb8)) ?
                  (wire114 ? reg119 : reg124) : wire112[(4'h8):(3'h4)]))));
              reg125 <= $signed($signed($signed($unsigned(wire114[(2'h2):(1'h1)]))));
              reg126 <= $signed(reg121);
            end
          else
            begin
              reg124 <= $signed(reg126);
              reg125 <= $unsigned((((7'h42) ?
                      reg122 : $signed({reg119, wire123})) ?
                  (-(wire116[(1'h0):(1'h0)] ?
                      wire117 : (wire114 ?
                          (7'h40) : reg119))) : ((~$unsigned(wire117)) ?
                      (&$unsigned(reg119)) : reg124)));
              reg126 <= wire114;
              reg127 <= $signed(reg126);
              reg128 <= (&($unsigned(wire113[(2'h3):(1'h1)]) ?
                  (+(-wire112)) : $signed($unsigned({reg119}))));
            end
          reg129 <= $unsigned(reg128);
          reg130 <= ((!(~reg126[(3'h7):(3'h5)])) ?
              (~&{wire120[(3'h5):(3'h4)],
                  $unsigned($unsigned(wire114))}) : reg124);
        end
      reg131 <= ((8'hb5) ?
          {wire117[(2'h2):(1'h0)],
              (((wire113 >= wire117) * reg125) ?
                  (^~{reg130}) : $unsigned($signed((8'ha9))))} : $unsigned(wire113[(2'h3):(2'h3)]));
      reg132 <= reg131[(3'h5):(2'h2)];
      reg133 <= $signed((+wire123[(2'h2):(2'h2)]));
      if (wire116[(4'h8):(4'h8)])
        begin
          reg134 <= (wire116 >= (^(8'hb2)));
        end
      else
        begin
          if (reg131)
            begin
              reg134 <= reg128;
              reg135 <= reg119;
              reg136 <= ($signed($unsigned($signed(reg125[(3'h6):(1'h1)]))) ^~ (reg134[(1'h1):(1'h0)] && $signed($unsigned(wire116[(3'h7):(3'h7)]))));
            end
          else
            begin
              reg134 <= (!((!$signed((reg127 < wire123))) == ((!reg127[(4'hf):(4'h9)]) ?
                  reg129 : wire115[(4'hc):(4'h8)])));
              reg135 <= $unsigned((~^((reg135[(3'h7):(3'h4)] ?
                  reg130[(3'h4):(2'h3)] : (~reg131)) != (~|$unsigned(wire112)))));
            end
          reg137 <= reg130;
          reg138 <= reg125;
          reg139 <= ((($signed(reg127[(4'hb):(2'h2)]) <<< $signed((&reg138))) * (reg124[(3'h6):(2'h2)] ?
                  (reg128 ~^ {(8'ha0), wire113}) : reg137[(3'h5):(2'h3)])) ?
              $unsigned(wire113[(4'hc):(2'h3)]) : ((wire114[(1'h0):(1'h0)] ?
                      {(reg131 << wire112)} : $unsigned((wire114 ?
                          reg130 : reg129))) ?
                  ($unsigned(reg136[(1'h1):(1'h0)]) ^~ $unsigned(reg133[(3'h7):(2'h2)])) : $unsigned({(~wire120),
                      wire113[(3'h5):(1'h0)]})));
          reg140 <= (((reg133[(2'h3):(1'h1)] <<< reg119) || (!$signed(wire113[(3'h7):(3'h4)]))) & {reg124[(1'h0):(1'h0)],
              $signed($signed($signed(wire113)))});
        end
    end
  assign wire141 = ({wire112} + (wire118[(1'h1):(1'h0)] ~^ reg130[(3'h4):(2'h2)]));
  assign wire142 = {reg128[(1'h0):(1'h0)], {((~|(&(8'ha0))) << (-(~^reg136)))}};
  assign wire143 = ((~wire120) ?
                       $unsigned((wire142[(4'he):(2'h3)] ?
                           wire115[(1'h1):(1'h0)] : wire141)) : {(~^(^~wire141))});
  assign wire144 = reg131;
  assign wire145 = (8'hb2);
  assign wire146 = $unsigned({(|(^reg137[(2'h2):(2'h2)])), wire120});
  always
    @(posedge clk) begin
      if ($unsigned($signed((+wire120[(4'h9):(4'h8)]))))
        begin
          reg147 <= (reg121 | {(~|($unsigned(wire123) ?
                  $unsigned(wire145) : $unsigned((8'haa))))});
          reg148 <= (wire144[(4'h8):(1'h1)] > ((-(+$unsigned((8'hba)))) ?
              {$signed(wire116[(1'h1):(1'h1)]), (^(~^(8'hb0)))} : (({(8'ha7),
                      (8'hb5)} ?
                  $unsigned(reg129) : $unsigned(reg127)) <= $signed((wire144 ?
                  wire116 : reg121)))));
          reg149 <= ($signed($unsigned((+(reg137 ? (8'haf) : reg148)))) ?
              $signed({((reg135 && reg137) > ((8'ha9) <= wire142)),
                  (~&(8'hae))}) : reg139);
          if ($signed(reg126[(1'h0):(1'h0)]))
            begin
              reg150 <= ((8'hbc) * $unsigned($unsigned($unsigned((~&(8'hac))))));
              reg151 <= $unsigned({$unsigned(reg136[(1'h0):(1'h0)])});
              reg152 <= (((-(8'ha1)) ? (8'ha0) : wire117) ?
                  $signed(reg138[(3'h6):(2'h2)]) : (~^($signed(((8'ha0) ?
                          reg133 : wire120)) ?
                      wire118[(1'h1):(1'h1)] : reg140[(4'ha):(2'h2)])));
              reg153 <= wire115;
              reg154 <= reg140[(3'h7):(3'h6)];
            end
          else
            begin
              reg150 <= $unsigned((8'ha0));
              reg151 <= {reg148, wire118[(3'h4):(2'h2)]};
              reg152 <= ((-(-wire141[(4'h9):(2'h3)])) ?
                  wire117 : (~((7'h43) ?
                      ($unsigned(reg137) - reg135[(4'hd):(1'h0)]) : ($unsigned((8'ha2)) ?
                          $unsigned(reg147) : (~|reg132)))));
              reg153 <= (8'ha2);
              reg154 <= (wire117[(4'h9):(1'h1)] <= $unsigned(wire144));
            end
          if ({(^$signed(($signed(reg131) ?
                  reg132[(4'he):(4'ha)] : (wire117 >> wire113))))})
            begin
              reg155 <= ($unsigned(wire146[(1'h1):(1'h0)]) ?
                  $signed((8'h9f)) : $signed((~|$signed(wire143[(2'h2):(1'h1)]))));
              reg156 <= (~^$signed(reg151[(1'h0):(1'h0)]));
              reg157 <= reg156;
            end
          else
            begin
              reg155 <= {wire146[(2'h2):(2'h2)],
                  ((reg119[(3'h6):(3'h6)] <<< $unsigned((reg153 ?
                          (7'h43) : (8'ha3)))) ?
                      (~^(|wire114[(2'h2):(1'h1)])) : (wire143[(1'h0):(1'h0)] <= (((8'hb6) ?
                              wire116 : reg126) ?
                          $signed(reg135) : $signed(wire142))))};
              reg156 <= (~|(|(~|reg127[(1'h1):(1'h1)])));
              reg157 <= ((reg131[(3'h5):(3'h5)] - {reg136[(3'h5):(1'h1)],
                  ($signed(wire117) && (^~reg130))}) < reg131[(4'h8):(1'h1)]);
              reg158 <= (($signed($signed({reg119})) - $signed($signed(reg122))) < $unsigned({reg132,
                  ($signed((8'ha1)) ? reg137[(2'h2):(1'h0)] : (8'hb4))}));
            end
        end
      else
        begin
          reg147 <= $signed(reg140[(4'ha):(1'h1)]);
          reg148 <= (wire123 * {wire142, (~reg134[(2'h2):(1'h0)])});
        end
      reg159 <= reg153[(2'h2):(2'h2)];
    end
  assign wire160 = $signed($unsigned($unsigned(((reg138 & (8'h9e)) ?
                       (reg134 < wire146) : {(8'h9f), (8'ha8)}))));
endmodule

module module78  (y, clk, wire82, wire81, wire80, wire79);
  output wire [(32'hcc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire82;
  input wire signed [(5'h15):(1'h0)] wire81;
  input wire [(3'h6):(1'h0)] wire80;
  input wire [(4'h8):(1'h0)] wire79;
  wire signed [(4'h9):(1'h0)] wire98;
  wire [(5'h10):(1'h0)] wire97;
  wire signed [(2'h3):(1'h0)] wire96;
  wire signed [(4'hb):(1'h0)] wire95;
  wire [(4'h8):(1'h0)] wire91;
  wire [(3'h4):(1'h0)] wire90;
  wire [(4'hb):(1'h0)] wire89;
  wire [(4'h9):(1'h0)] wire88;
  wire signed [(4'hb):(1'h0)] wire84;
  wire [(4'hb):(1'h0)] wire83;
  reg [(2'h2):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg100 = (1'h0);
  reg [(3'h4):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg94 = (1'h0);
  reg [(4'ha):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg92 = (1'h0);
  reg [(4'h8):(1'h0)] reg87 = (1'h0);
  reg [(5'h12):(1'h0)] reg86 = (1'h0);
  reg [(5'h15):(1'h0)] reg85 = (1'h0);
  assign y = {wire98,
                 wire97,
                 wire96,
                 wire95,
                 wire91,
                 wire90,
                 wire89,
                 wire88,
                 wire84,
                 wire83,
                 reg101,
                 reg100,
                 reg99,
                 reg94,
                 reg93,
                 reg92,
                 reg87,
                 reg86,
                 reg85,
                 (1'h0)};
  assign wire83 = wire80[(3'h5):(3'h5)];
  assign wire84 = (((~$signed((|wire82))) ?
                          (wire79[(4'h8):(2'h2)] ~^ ($signed(wire80) ?
                              $signed(wire82) : $signed(wire81))) : ((((8'hb1) > (8'hbc)) || $signed(wire82)) & $unsigned($unsigned((8'hbc))))) ?
                      (&($unsigned(wire82) ?
                          wire83[(1'h1):(1'h0)] : wire82[(1'h0):(1'h0)])) : wire81[(4'ha):(4'h9)]);
  always
    @(posedge clk) begin
      reg85 <= $signed(wire79[(3'h6):(2'h2)]);
      reg86 <= wire82;
      reg87 <= $signed({wire80[(2'h3):(2'h3)],
          (-(wire81 ? wire84[(1'h0):(1'h0)] : wire82[(1'h1):(1'h0)]))});
    end
  assign wire88 = (7'h41);
  assign wire89 = {(^~wire80)};
  assign wire90 = reg87;
  assign wire91 = ($signed($signed((~^wire83[(2'h3):(1'h1)]))) ?
                      (&$unsigned((wire90 | ((8'ha5) ?
                          reg87 : wire90)))) : (!({{wire84}} == (wire89[(3'h6):(2'h3)] - (wire83 ?
                          wire84 : wire90)))));
  always
    @(posedge clk) begin
      if ({(+$unsigned(reg85)),
          ($signed((~&((8'ha2) < wire83))) & $unsigned((wire82[(1'h0):(1'h0)] ?
              wire91[(1'h1):(1'h0)] : $signed(reg86))))})
        begin
          reg92 <= (~{((wire79 ^~ $signed(reg86)) && wire81)});
          reg93 <= ((^{$signed((wire88 | wire81))}) * (!$unsigned($unsigned($unsigned(wire80)))));
          reg94 <= wire81;
        end
      else
        begin
          reg92 <= $signed(wire79);
          reg93 <= reg93;
        end
    end
  assign wire95 = (+(~&wire80[(3'h4):(1'h0)]));
  assign wire96 = reg92[(4'hc):(1'h1)];
  assign wire97 = $signed($unsigned(reg93[(3'h6):(3'h4)]));
  assign wire98 = {(&wire84[(3'h5):(3'h4)]),
                      ((7'h43) ?
                          wire80[(1'h1):(1'h0)] : $signed((((8'ha6) << wire82) != $unsigned(reg86))))};
  always
    @(posedge clk) begin
      reg99 <= {$signed({(+wire95[(1'h1):(1'h1)]), (reg94 || wire81)}),
          (wire81[(4'he):(3'h5)] ?
              (~&($unsigned(wire79) ?
                  (wire84 || wire91) : ((8'hb4) ?
                      wire80 : wire82))) : (+{wire90[(1'h1):(1'h1)],
                  $signed((8'hac))}))};
      reg100 <= wire95;
      reg101 <= $unsigned((^~(&$unsigned($signed(wire96)))));
    end
endmodule

module module23
#(parameter param73 = (~|(((((7'h40) ? (8'haf) : (8'ha3)) != ((8'h9c) ? (8'ha9) : (8'haa))) ? (|(^(8'hb5))) : {((8'ha2) > (8'ha4)), ((8'ha2) - (8'had))}) ? ((((8'hb8) ? (8'ha0) : (8'hb0)) * {(7'h42), (8'had)}) && ((~|(8'hb5)) + ((8'hb3) ? (8'hbb) : (7'h43)))) : (~&(^~((8'ha3) ? (8'hb4) : (8'ha3)))))))
(y, clk, wire27, wire26, wire25, wire24);
  output wire [(32'h251):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire27;
  input wire [(2'h2):(1'h0)] wire26;
  input wire [(3'h4):(1'h0)] wire25;
  input wire [(3'h5):(1'h0)] wire24;
  wire [(4'hb):(1'h0)] wire72;
  wire signed [(4'he):(1'h0)] wire71;
  wire signed [(4'hb):(1'h0)] wire62;
  wire signed [(2'h3):(1'h0)] wire61;
  wire signed [(5'h13):(1'h0)] wire60;
  wire [(4'ha):(1'h0)] wire59;
  wire [(3'h7):(1'h0)] wire58;
  wire signed [(5'h11):(1'h0)] wire57;
  wire [(4'hd):(1'h0)] wire56;
  wire [(4'he):(1'h0)] wire55;
  wire [(5'h13):(1'h0)] wire54;
  wire signed [(5'h10):(1'h0)] wire53;
  wire signed [(4'hb):(1'h0)] wire52;
  wire signed [(5'h12):(1'h0)] wire51;
  wire signed [(5'h14):(1'h0)] wire50;
  wire [(4'h9):(1'h0)] wire43;
  wire [(4'hf):(1'h0)] wire42;
  wire signed [(5'h12):(1'h0)] wire41;
  wire signed [(4'hf):(1'h0)] wire40;
  reg signed [(5'h12):(1'h0)] reg70 = (1'h0);
  reg [(5'h10):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg68 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg67 = (1'h0);
  reg [(4'ha):(1'h0)] reg66 = (1'h0);
  reg [(3'h6):(1'h0)] reg65 = (1'h0);
  reg [(4'he):(1'h0)] reg64 = (1'h0);
  reg [(4'hb):(1'h0)] reg63 = (1'h0);
  reg [(3'h7):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg48 = (1'h0);
  reg [(4'ha):(1'h0)] reg47 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg46 = (1'h0);
  reg [(4'hb):(1'h0)] reg45 = (1'h0);
  reg [(5'h15):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg39 = (1'h0);
  reg [(5'h11):(1'h0)] reg38 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg37 = (1'h0);
  reg [(5'h13):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg34 = (1'h0);
  reg signed [(4'he):(1'h0)] reg33 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg31 = (1'h0);
  reg [(5'h12):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg29 = (1'h0);
  reg [(4'hc):(1'h0)] reg28 = (1'h0);
  assign y = {wire72,
                 wire71,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire43,
                 wire42,
                 wire41,
                 wire40,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(wire24)))
        begin
          reg28 <= wire27[(1'h1):(1'h0)];
          if (reg28)
            begin
              reg29 <= wire25[(3'h4):(1'h1)];
              reg30 <= $signed({$unsigned(wire25)});
              reg31 <= $unsigned(((-$signed((^wire25))) ?
                  ({$unsigned(wire24),
                      reg29} - $unsigned(reg30)) : ($unsigned((^(8'ha0))) == wire25)));
              reg32 <= $unsigned(((^~(wire24 <<< $unsigned(reg28))) ?
                  (~|$unsigned($unsigned(reg29))) : {wire24}));
              reg33 <= reg31;
            end
          else
            begin
              reg29 <= (^$signed((~|reg28[(2'h3):(2'h3)])));
              reg30 <= $signed((+wire25));
              reg31 <= (8'ha5);
              reg32 <= $signed(((wire25 && $unsigned((8'hac))) > reg30[(3'h6):(3'h5)]));
              reg33 <= (-(({$unsigned(reg29), $unsigned(wire25)} ?
                      ((reg30 + reg28) ^ $signed(reg29)) : reg30) ?
                  reg31[(5'h11):(4'hf)] : {(((8'had) * wire26) ?
                          wire27 : $unsigned(reg32)),
                      {$unsigned(reg32)}}));
            end
          reg34 <= wire26[(2'h2):(1'h0)];
          if ((reg28 * {(~&$signed(reg28[(1'h0):(1'h0)])),
              $unsigned($signed((^reg29)))}))
            begin
              reg35 <= $signed(reg31);
              reg36 <= $unsigned(reg28);
              reg37 <= (~|$signed(wire25));
            end
          else
            begin
              reg35 <= reg29[(5'h11):(4'hf)];
              reg36 <= (wire27[(3'h7):(3'h5)] ?
                  ((^~reg31[(4'hc):(4'hb)]) == ($unsigned((reg35 == reg35)) ?
                      wire26[(2'h2):(2'h2)] : (^(reg37 >>> wire25)))) : (~|(8'ha1)));
              reg37 <= {($unsigned((|(wire26 ? reg36 : (8'hbb)))) ?
                      $signed(((reg30 ? reg30 : reg29) ^~ (8'ha6))) : reg34)};
              reg38 <= (7'h42);
            end
        end
      else
        begin
          reg28 <= reg34[(4'ha):(4'h8)];
          reg29 <= $signed(wire27[(2'h2):(2'h2)]);
          reg30 <= (({((reg36 ? reg32 : (8'hba)) ? {wire27} : (reg29 ^ wire24)),
                  $signed((|reg33))} ?
              (^~(!$unsigned(reg29))) : reg36[(3'h5):(3'h4)]) >> ({(!$unsigned(reg28)),
                  reg29[(5'h13):(3'h7)]} ?
              $signed($signed((reg37 ? reg30 : reg38))) : ((8'hb6) ?
                  wire24[(1'h1):(1'h1)] : (|(-reg35)))));
          reg31 <= $signed(reg32);
        end
      reg39 <= (((8'ha7) >>> $signed(((reg31 * (8'ha9)) ~^ reg34[(4'hc):(4'hc)]))) ?
          $unsigned(((^reg38[(3'h7):(2'h3)]) | reg32)) : (+$signed($signed($signed(wire27)))));
    end
  assign wire40 = (&(~&$unsigned(reg33[(4'h8):(3'h5)])));
  assign wire41 = ((($unsigned(wire27) || reg32[(1'h0):(1'h0)]) ?
                      ($unsigned((wire25 > (8'ha7))) << ((reg32 ^~ wire40) && reg33)) : reg31[(3'h6):(1'h1)]) && ({reg31,
                      (+{reg35, reg36})} < (~$signed(wire25[(3'h4):(1'h1)]))));
  assign wire42 = (+wire27);
  assign wire43 = (~^({{$signed(reg30)}} ?
                      $signed((~|$unsigned(wire41))) : wire41[(4'ha):(4'h9)]));
  always
    @(posedge clk) begin
      if (reg38)
        begin
          reg44 <= ((~^$signed(({wire27} | {wire42}))) ?
              (($unsigned({reg38, (8'ha3)}) ^~ wire41[(3'h7):(2'h3)]) ?
                  $signed((~$signed(reg39))) : $signed({(wire25 ?
                          reg39 : (8'ha7)),
                      reg39})) : ((8'h9c) & (~&$unsigned((reg31 != (7'h43))))));
          reg45 <= reg35;
          reg46 <= reg37[(1'h1):(1'h0)];
          if (($signed($signed((+$signed(reg36)))) <<< {(reg28[(4'h8):(4'h8)] ?
                  $unsigned((wire40 >= reg36)) : (8'ha2))}))
            begin
              reg47 <= {(reg44[(5'h13):(4'he)] ?
                      $signed({reg37}) : reg33[(4'h8):(4'h8)])};
              reg48 <= ($signed((($signed((8'hba)) >> $unsigned(reg31)) >= $unsigned((reg45 ?
                      wire43 : (8'hab))))) ?
                  ($unsigned((~&(8'h9f))) ?
                      ($signed({reg38, wire27}) ?
                          ($unsigned(reg44) * ((8'hbd) ?
                              wire43 : wire41)) : wire25) : ((^reg45) * $signed(wire27))) : wire24[(1'h1):(1'h1)]);
              reg49 <= ($unsigned((+reg46[(3'h5):(2'h3)])) ?
                  wire26[(1'h0):(1'h0)] : reg28);
            end
          else
            begin
              reg47 <= (reg46[(3'h6):(1'h1)] ?
                  ((~|reg47) ?
                      (~|reg44[(3'h6):(3'h6)]) : ((~&(^(8'hbc))) ?
                          $signed($unsigned(reg32)) : $signed((^reg44)))) : reg45);
              reg48 <= {(^($signed(wire26) ?
                      ({reg46} ?
                          (~^(8'hae)) : $signed(wire26)) : $signed({reg39}))),
                  $signed($signed({((7'h43) ? reg34 : wire43)}))};
            end
        end
      else
        begin
          if ($signed((^(~$signed(reg37[(1'h1):(1'h0)])))))
            begin
              reg44 <= ((($signed(reg46) ?
                      $unsigned(reg28[(4'h9):(2'h2)]) : $unsigned((reg30 ^~ wire42))) >>> (^~(reg28 ~^ reg29))) ?
                  $unsigned(($unsigned((reg33 ? (8'hb1) : reg39)) ?
                      $signed($signed(reg33)) : {$unsigned(reg29)})) : $unsigned({$unsigned(((7'h43) ?
                          reg44 : reg28)),
                      reg28[(2'h3):(2'h2)]}));
              reg45 <= {wire40[(1'h0):(1'h0)],
                  ({$signed(reg45), reg33[(1'h1):(1'h1)]} <<< (!reg37))};
              reg46 <= (^~reg36);
              reg47 <= reg31[(4'ha):(1'h1)];
              reg48 <= ({reg32, wire43[(1'h0):(1'h0)]} ?
                  {$unsigned($signed(wire24)),
                      $unsigned(((reg31 * (8'hbf)) && wire42[(4'hb):(1'h0)]))} : ({{$unsigned(reg28),
                          (|wire43)}} <= wire26));
            end
          else
            begin
              reg44 <= ((($unsigned(wire24) ^ reg36[(3'h7):(1'h0)]) >= (8'ha1)) ?
                  wire26[(2'h2):(1'h0)] : reg48[(3'h5):(2'h3)]);
              reg45 <= (&((7'h43) << (reg45[(2'h3):(2'h2)] <<< $unsigned(wire41[(4'hc):(4'hb)]))));
              reg46 <= (^~reg29[(5'h12):(4'ha)]);
              reg47 <= ($unsigned({(&(reg29 ? reg33 : reg35)),
                  ({wire24, reg28} ^~ (wire43 ?
                      (8'hbe) : reg38))}) && (({$unsigned(reg46)} ?
                      (^(reg29 ? reg46 : (8'hba))) : (~|(-reg47))) ?
                  (($unsigned(reg37) << (wire43 ?
                      wire40 : wire41)) <= $unsigned((reg38 & wire26))) : $signed(wire40)));
              reg48 <= {(^$unsigned($signed($unsigned(reg35)))),
                  ((8'ha4) ? reg35 : $signed((reg45 != $unsigned(reg47))))};
            end
        end
    end
  assign wire50 = reg48[(2'h3):(1'h0)];
  assign wire51 = {(|wire41[(3'h4):(2'h2)])};
  assign wire52 = (~|wire51[(3'h7):(3'h5)]);
  assign wire53 = $unsigned((~|reg47));
  assign wire54 = ((^~(~|$signed($unsigned(reg44)))) ?
                      wire25[(3'h4):(1'h0)] : (|reg49[(1'h1):(1'h1)]));
  assign wire55 = (reg35 ?
                      $signed((reg39 ?
                          (^{reg49}) : reg35[(3'h5):(3'h5)])) : ((~^wire25) ?
                          wire52[(2'h3):(1'h0)] : {wire52[(3'h7):(2'h2)]}));
  assign wire56 = ($signed({(-(reg38 < (8'hb0))), (^~{reg35, reg45})}) ?
                      {$signed((wire40[(1'h1):(1'h0)] ?
                              $signed(reg29) : $signed(reg36)))} : (^(-(^~$signed(reg45)))));
  assign wire57 = ((^~(!reg39[(3'h6):(3'h5)])) ?
                      {$unsigned(reg29[(4'ha):(3'h6)])} : ({reg44[(2'h3):(2'h3)],
                              {reg33}} ?
                          wire24 : $signed(wire50)));
  assign wire58 = $unsigned((+((wire55 == wire40[(3'h6):(1'h0)]) + ((wire50 ?
                          wire25 : wire53) ?
                      (reg31 == reg47) : wire56[(2'h2):(2'h2)]))));
  assign wire59 = wire25[(1'h1):(1'h1)];
  assign wire60 = $signed({(reg44 >> ($signed(reg32) >>> (wire43 * reg30))),
                      wire50[(3'h5):(3'h4)]});
  assign wire61 = $signed(((-(((8'hb7) ~^ wire56) * $signed(wire43))) && reg34[(1'h1):(1'h0)]));
  assign wire62 = $signed((8'hbc));
  always
    @(posedge clk) begin
      if ((((reg38[(4'h9):(4'h8)] ?
                  $unsigned(reg33[(3'h5):(2'h3)]) : ($signed(reg33) ?
                      (wire54 ? reg31 : reg33) : reg38[(1'h0):(1'h0)])) ?
              $unsigned((wire52 || (-(8'hbf)))) : $signed($signed((reg37 ?
                  wire61 : wire57)))) ?
          reg30 : (&((^~$signed(wire53)) != ({reg39, reg36} != (wire62 ?
              wire54 : (8'hb0)))))))
        begin
          reg63 <= $unsigned((|$signed($signed((-wire57)))));
          reg64 <= $signed((reg38[(1'h0):(1'h0)] < $signed($unsigned((~|reg47)))));
          reg65 <= (^($unsigned(((!wire59) >>> {reg28,
              reg45})) ^~ ($signed({(8'hbd)}) ?
              $signed((wire56 != wire54)) : $signed((wire41 ?
                  reg38 : reg32)))));
          if ($unsigned($unsigned(wire50)))
            begin
              reg66 <= $signed((((^((8'h9f) >= wire56)) + (wire60[(2'h3):(1'h1)] ?
                      reg30[(1'h0):(1'h0)] : ((7'h42) && (8'ha5)))) ?
                  reg49 : wire57));
              reg67 <= $unsigned($unsigned(reg64[(4'hd):(4'hb)]));
            end
          else
            begin
              reg66 <= wire55[(2'h3):(1'h1)];
              reg67 <= ($unsigned(reg31[(4'he):(4'h8)]) ?
                  wire24[(1'h0):(1'h0)] : (^reg64));
            end
        end
      else
        begin
          reg63 <= $signed((reg39 < reg65));
          reg64 <= wire58;
          if ((($unsigned(reg29[(4'he):(4'hd)]) ?
              {{reg66}} : ($unsigned(reg29[(5'h11):(4'hd)]) * $unsigned(((7'h44) < wire53)))) | (8'hb6)))
            begin
              reg65 <= (~$unsigned((wire52[(2'h2):(1'h1)] ^~ $signed((reg64 ?
                  wire41 : wire59)))));
              reg66 <= (+($signed((reg49[(3'h5):(2'h2)] ?
                  (reg47 ?
                      reg47 : wire40) : wire52[(1'h1):(1'h0)])) < ($signed($unsigned(reg28)) ?
                  (|reg48) : {(reg31 ? reg29 : (8'hbb))})));
              reg67 <= $signed($signed((!$unsigned($unsigned((8'had))))));
            end
          else
            begin
              reg65 <= (((&wire42[(3'h5):(1'h1)]) ?
                      reg45[(4'h9):(4'h8)] : {{$signed(reg46)},
                          $signed($signed(wire58))}) ?
                  $unsigned($signed((reg32 ?
                      reg66 : (~^wire56)))) : (~|$unsigned({reg49[(2'h2):(1'h1)],
                      reg46[(4'ha):(4'h8)]})));
              reg66 <= wire50[(2'h2):(1'h1)];
            end
        end
      reg68 <= (8'ha6);
      reg69 <= (-$signed((wire54 ?
          ((reg64 + reg36) > $signed(reg63)) : reg35[(3'h7):(3'h5)])));
      reg70 <= {reg44};
    end
  assign wire71 = reg39;
  assign wire72 = wire58[(2'h2):(1'h0)];
endmodule
